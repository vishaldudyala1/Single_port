vas,fm
