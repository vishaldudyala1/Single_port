gkhajk
